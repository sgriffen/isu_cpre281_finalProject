module Input_Logic_TLC_Mk3 (en, w, y, X);
	
	input en;
	input [1:0]w;
	input [3:0]y;
	output [3:0]X;
	
	reg [3:0]X;
	
	always @(en or w or y)
	begin
		case({en, w, y})
			
			//Count up (Add car)
			7'b 1010000: X = 4'b 0001; //A
			7'b 1010001: X = 4'b 0010; //B
			7'b 1010010: X = 4'b 0011; //C
			7'b 1010011: X = 4'b 0100; //D
			7'b 1010100: X = 4'b 0101; //E
			7'b 1010101: X = 4'b 0110; //F
			7'b 1010110: X = 4'b 0111; //G
			7'b 1010111: X = 4'b 1000; //H
			7'b 1011000: X = 4'b 1001; //I
			7'b 1011001: X = 4'b 1010; //J
			7'b 1011010: X = 4'b 1011; //K
			7'b 1011011: X = 4'b 1100; //L
			7'b 1011100: X = 4'b 1101; //M
			7'b 1011101: X = 4'b 1110; //N
			7'b 1011110: X = 4'b 1111; //O
			7'b 1011111: X = 4'b 1111; //P
			
			//Count down (Green light)
			7'b 1100000: X = 4'b 0000; //A
			7'b 1100001: X = 4'b 0000; //B
			7'b 1100010: X = 4'b 0001; //C
			7'b 1100011: X = 4'b 0010; //D
			7'b 1100100: X = 4'b 0011; //E
			7'b 1100101: X = 4'b 0100; //F
			7'b 1100110: X = 4'b 0101; //G
			7'b 1100111: X = 4'b 0110; //H
			7'b 1101000: X = 4'b 0111; //I
			7'b 1101001: X = 4'b 1000; //J
			7'b 1101010: X = 4'b 1001; //K
			7'b 1101011: X = 4'b 1010; //L
			7'b 1101100: X = 4'b 1011; //M
			7'b 1101101: X = 4'b 1100; //N
			7'b 1101110: X = 4'b 1101; //O
			7'b 1101111: X = 4'b 1110; //P
			
			//Default Cases
			7'b 0000000: X = 4'b 0000;
			7'b 0000001: X = 4'b 0001;
			7'b 0000010: X = 4'b 0010;
			7'b 0000011: X = 4'b 0011;
			7'b 0000100: X = 4'b 0100;
			7'b 0000101: X = 4'b 0101;
			7'b 0000110: X = 4'b 0110;
			7'b 0000111: X = 4'b 0111;
			7'b 0001000: X = 4'b 1000;
			7'b 0001001: X = 4'b 1001;
			7'b 0001010: X = 4'b 1010;
			7'b 0001011: X = 4'b 1011;
			7'b 0001100: X = 4'b 1100;
			7'b 0001101: X = 4'b 1101;
			7'b 0001110: X = 4'b 1110;
			7'b 0001111: X = 4'b 1111;
			
			7'b 0010000: X = 4'b 0000;
			7'b 0010001: X = 4'b 0001;
			7'b 0010010: X = 4'b 0010;
			7'b 0000011: X = 4'b 0011;
			7'b 0010100: X = 4'b 0100;
			7'b 0010101: X = 4'b 0101;
			7'b 0010110: X = 4'b 0110;
			7'b 0010111: X = 4'b 0111;
			7'b 0011000: X = 4'b 1000;
			7'b 0011001: X = 4'b 1001;
			7'b 0011010: X = 4'b 1010;
			7'b 0011011: X = 4'b 1011;
			7'b 0011100: X = 4'b 1100;
			7'b 0011101: X = 4'b 1101;
			7'b 0011110: X = 4'b 1110;
			7'b 0011111: X = 4'b 1111;
			
			7'b 0100000: X = 4'b 0000;
			7'b 0100001: X = 4'b 0001;
			7'b 0100010: X = 4'b 0010;
			7'b 0100011: X = 4'b 0011;
			7'b 0100100: X = 4'b 0100;
			7'b 0100101: X = 4'b 0101;
			7'b 0100110: X = 4'b 0110;
			7'b 0100111: X = 4'b 0111;
			7'b 0101000: X = 4'b 1000;
			7'b 0101001: X = 4'b 1001;
			7'b 0101010: X = 4'b 1010;
			7'b 0101011: X = 4'b 1011;
			7'b 0101100: X = 4'b 1100;
			7'b 0101101: X = 4'b 1101;
			7'b 0101110: X = 4'b 1110;
			7'b 0101111: X = 4'b 1111;
			
			7'b 0110000: X = 4'b 0000;
			7'b 0110001: X = 4'b 0001;
			7'b 0110010: X = 4'b 0010;
			7'b 0110011: X = 4'b 0011;
			7'b 0110100: X = 4'b 0100;
			7'b 0110101: X = 4'b 0101;
			7'b 0110110: X = 4'b 0110;
			7'b 0110111: X = 4'b 0111;
			7'b 0111000: X = 4'b 1000;
			7'b 0111001: X = 4'b 1001;
			7'b 0111010: X = 4'b 1010;
			7'b 0111011: X = 4'b 1011;
			7'b 0111100: X = 4'b 1100;
			7'b 0111101: X = 4'b 1101;
			7'b 0111110: X = 4'b 1110;
			7'b 0111111: X = 4'b 1111;
		
			7'b 1000000: X = 4'b 0000;
			7'b 1000001: X = 4'b 0001;
			7'b 1000010: X = 4'b 0010;
			7'b 1000011: X = 4'b 0011;
			7'b 1000100: X = 4'b 0100;
			7'b 1000101: X = 4'b 0101;
			7'b 1000110: X = 4'b 0110;
			7'b 1000111: X = 4'b 0111;
			7'b 1001000: X = 4'b 1000;
			7'b 1001001: X = 4'b 1001;
			7'b 1001010: X = 4'b 1010;
			7'b 1001011: X = 4'b 1011;
			7'b 1001100: X = 4'b 1100;
			7'b 1001101: X = 4'b 1101;
			7'b 1001110: X = 4'b 1110;
			7'b 1001111: X = 4'b 1111;
		
			7'b 1110000: X = 4'b 0000;
			7'b 1110001: X = 4'b 0001;
			7'b 1110010: X = 4'b 0010;
			7'b 1110011: X = 4'b 0011;
			7'b 1110100: X = 4'b 0100;
			7'b 1110101: X = 4'b 0101;
			7'b 1110110: X = 4'b 0110;
			7'b 1110111: X = 4'b 0111;
			7'b 1111000: X = 4'b 1000;
			7'b 1111001: X = 4'b 1001;
			7'b 1111010: X = 4'b 1010;
			7'b 1111011: X = 4'b 1011;
			7'b 1111100: X = 4'b 1100;
			7'b 1111101: X = 4'b 1101;
			7'b 1111110: X = 4'b 1110;
			7'b 1111111: X = 4'b 1111;
			
		endcase
	end
endmodule