module Input_Logic (w, y, X);

	input w;
	input [3:0]y;
	output [3:0]X;
		
	assign X[3] = (y[3] & y[2])|(y[3] & y[1])|(y[3] & y[0])|(w & y[3])|(w & y[2] & y[1] & y[0]);
	assign X[2] = (y[2] & ~y[1] & y[0]) | (y[2] & y[1] & ~y[0]) | (~w & y[2] & y[1]) | (w & y[2] & ~y[1]) | (w & y[3] & y[1] & y[0]) | (w & ~y[2] & y[1] & y[0]) | (~w & y[3] & ~y[2] & ~y[1] & ~y[0]);
	assign X[1] = (~w & y[1] & y[0]) | (~w & y[2] & ~y[1] & ~y[0]) | (~w & y[3] & ~y[1] & ~y[0]) | (w & y[1] & ~y[0]) | (w & ~y[1] & y[0]) | (w & y[3] & y[2] & y[0]);
	assign X[0] = (y[1] & ~y[0]) | (y[3] & ~y[0]) | (y[2] & ~y[0]) | (w & ~y[3] & ~y[0]) | (w & y[3] & y[2] & y[1]);
	
endmodule