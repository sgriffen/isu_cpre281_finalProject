module Input_Logic_TLC_Mk2 (w, y, X);

	input [1:0]w;
	input [3:0]y;
	output [3:0]X;
	
	reg [3:0]X;
	
	always @(w or y)
	begin
		case(w)
		
			2'b 01: X = {(y[3] & y[2])|(y[3] & y[1])|(y[3] & y[0])|(w[0] & y[3])|(w[0] & y[2] & y[1] & y[0]),
							 (y[2] & ~y[1] & y[0]) | (y[2] & y[1] & ~y[0]) | (~w[0] & y[2] & y[1]) | (w[0] & y[2] & ~y[1]) | (w[0] & y[3] & y[1] & y[0]) | (w[0] & ~y[2] & y[1] & y[0]) | (~w[0] & y[3] & ~y[2] & ~y[1] & ~y[0]),
							  (~w[0] & y[1] & y[0]) | (~w[0] & y[2] & ~y[1] & ~y[0]) | (~w[0] & y[3] & ~y[1] & ~y[0]) | (w[0] & y[1] & ~y[0]) | (w[0] & ~y[1] & y[0]) | (w[0] & y[3] & y[2] & y[0]),
							  (y[1] & ~y[0]) | (y[3] & ~y[0]) | (y[2] & ~y[0]) | (w[0] & ~y[3] & ~y[0]) | (w[0] & y[3] & y[2] & y[1])};
			2'b 10: X = {(y[3] & y[2])|(y[3] & y[1])|(y[3] & y[0])|(w[0] & y[3])|(w[0] & y[2] & y[1] & y[0]),
							 (y[2] & ~y[1] & y[0]) | (y[2] & y[1] & ~y[0]) | (~w[0] & y[2] & y[1]) | (w[0] & y[2] & ~y[1]) | (w[0] & y[3] & y[1] & y[0]) | (w[0] & ~y[2] & y[1] & y[0]) | (~w[0] & y[3] & ~y[2] & ~y[1] & ~y[0]),
							  (~w[0] & y[1] & y[0]) | (~w[0] & y[2] & ~y[1] & ~y[0]) | (~w[0] & y[3] & ~y[1] & ~y[0]) | (w[0] & y[1] & ~y[0]) | (w[0] & ~y[1] & y[0]) | (w[0] & y[3] & y[2] & y[0]),
							  (y[1] & ~y[0]) | (y[3] & ~y[0]) | (y[2] & ~y[0]) | (w[0] & ~y[3] & ~y[0]) | (w[0] & y[3] & y[2] & y[1])};
			default: X = X;
		endcase
	end
endmodule